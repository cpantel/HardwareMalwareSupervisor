module counter(
   input CLK,
   input reset,
   input enable,
   input step,
   input fast,
   output reg [31:0] count,
   output reg running,
   output humanClock
);

initial count   = 0;

assign humanClock = fast ? count[24] : count[27];

always @(posedge CLK) 
begin
  if (reset) 
  begin
    count   <= 0;
  end 
  else if (enable) 
  begin
    count   <= count + 1;
  end
  else if (step) 
  begin
    count   <= count + 1;
  end
end
endmodule
