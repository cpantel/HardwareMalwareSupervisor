`timescale 1ns/1ps

module rom (
  input Clock,
  input reset,
  input [5:0] address,
  output reg [7:0] data
);
 
  reg [7:0]mem[0:47];

  always@(posedge Clock) begin
    case(address)
      16: data = 8'h90;  // nop
      17: data = 8'h90;  // nop  
      18: data = 8'h90;  // nop
      19: data = 8'h90;  // nop
      20: data = 8'h90;  // nop
      21: data = 8'h90;  // nop
      22: data = 8'h25;  // set   legal out
      23: data = 8'h40;  // svc
      24: data = 8'h2A;  // set
      25: data = 8'h40;  // svc
      26: data = 8'h2F;  // set
      27: data = 8'h40;  // svc
      28: data = 8'h25;  // set   failed out
      29: data = 8'h30;  // out
      30: data = 8'h2A;  // set
      31: data = 8'h30;  // out
      32: data = 8'h2F;  // set
      33: data = 8'h30;  // out
      34: data = 8'h20;  // set   troyan activation
      35: data = 8'h80;  // inc
      36: data = 8'h90;  // nop
      37: data = 8'h1F;  // jnz
      38: data = 8'h25;  // set   exploitation
      39: data = 8'h30;  // out   exploitation
      40: data = 8'h2A;  // set   exploitation
      41: data = 8'h30;  // out   exploitation
      42: data = 8'h2F;  // set   exploitation
      43: data = 8'h30;  // out   exploitation
      44: data = 8'h90;  // nop
      45: data = 8'h70;  // hlt
      46: data = 8'h30;  // out   svc
      47: data = 8'h00;  // ret
      default: data = 8'h00;
    endcase
    data =  mem[address];
  end
  
  
  always@(posedge reset)
   begin
   
    mem[0] = 8'h00;
    mem[1] = 8'h00;
    mem[2] = 8'h00;
    mem[3] = 8'h00;
    mem[4] = 8'h00;
    mem[5] = 8'h00;
    mem[6] = 8'h00;
    mem[7] = 8'h00;
    mem[8] = 8'h00;
    mem[9] = 8'h00;
    mem[10] = 8'h00;
    mem[11] = 8'h00;
    mem[12] = 8'h00;
    mem[13] = 8'h00;
    mem[14] = 8'h00;
    mem[15] = 8'h2e;
    mem[16] = 8'h90;
    mem[17] = 8'h90;
    mem[18] = 8'h90;
    mem[19] = 8'h90;
    mem[20] = 8'h90;
    mem[21] = 8'h90;
    mem[22] = 8'h25;
    mem[23] = 8'h40;
    mem[24] = 8'h2A;
    mem[25] = 8'h40;
    mem[26] = 8'h2F;
    mem[27] = 8'h40;
    mem[28] = 8'h25;
    mem[29] = 8'h30;
    mem[30] = 8'h2A;
    mem[31] = 8'h30;
    mem[32] = 8'h2F;
    mem[33] = 8'h30;
    mem[34] = 8'h20;
    mem[35] = 8'h80;
    mem[36] = 8'h90;
    mem[37] = 8'h1F;
    mem[38] = 8'h25;
    mem[39] = 8'h30;
    mem[40] = 8'h2A;
    mem[41] = 8'h30;
    mem[42] = 8'h2F;
    mem[43] = 8'h30;
    mem[44] = 8'h90;
    mem[45] = 8'h70;
    mem[46] = 8'h30;
    mem[47] = 8'h00;
  end
  
 
endmodule
