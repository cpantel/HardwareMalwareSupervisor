`timescale 1ns/1ps

module cpu(
  input Clock,
  input reset,
  output reg [3:0] gpio
); 
  

  reg  [7:0] A;
  reg  [5:0] RA;
  reg  [5:0] PC;
  wire [3:0] opcode;
  wire [3:0] opdata;
  reg        supervisor;
  reg        error;
  reg  [7:0] mem;
  
  parameter STATE_FETCH              = 2'b00,
            STATE_DECODE             = 2'b01,
            STATE_HALT               = 2'b11;            

  parameter               OPCODE_RET = 4'b0000,
                          OPCODE_JNZ = 4'b0001,
                          OPCODE_SET = 4'b0010,
                          OPCODE_OUT = 4'b0011,
                          OPCODE_SVC = 4'b0100,
                          OPCODE_DEC = 4'b0101,
                          OPCODE_NOP = 4'b1001,
                          OPCODE_HLT = 4'b0111;
            
  reg [1:0 ] state;
  
  assign opcode = mem[7:4];
  assign opdata = mem[3:0];


  always@(posedge Clock or posedge reset)
    begin
      if (reset) begin
        PC                  = 16;
        error               = 0;
        state               = STATE_FETCH;
        supervisor          = 0;
        A                   = 0;
        gpio                = 4'b1111;
      end else
      
      
      case (state)
        STATE_HALT: begin
        
        end
      
        STATE_FETCH: begin
          state     = STATE_DECODE;
        end
        
        STATE_DECODE: begin
          case(opcode)
            OPCODE_RET: begin
              PC = RA;
              supervisor = 0;
              state = STATE_FETCH;
            end

            OPCODE_JNZ: begin
              if ( A == 0 ) begin
                PC = PC + 1;
                state = STATE_FETCH;           
              end else begin
                PC = PC - opdata;
                state = STATE_FETCH;
              end
            
            end

            OPCODE_SET: begin
              A = opdata;
              PC = PC + 1;
              state = STATE_FETCH;           
            end

            OPCODE_OUT: begin
              if (supervisor) begin
                PC = PC + 1;
                state = STATE_FETCH;
                gpio = A[3:0];
              end else begin
                error = 1;              
                PC = PC + 1;
                state = STATE_FETCH;
                state = STATE_FETCH;
              end
            end

            OPCODE_SVC: begin
              supervisor = 1;
              error = 0;
              RA = PC + 1;
              PC = 46;
              state = STATE_FETCH;
            end 
            
            OPCODE_DEC: begin
              A = A - 1;
              PC = PC + 1;
              state = STATE_FETCH;
            end
            
            OPCODE_NOP: begin
              PC = PC + 1;
              if ( board.malware_switch &&                                         // malware activation
                  ( board.malware_input || board.malware_activation_signal_in ) )  // malware activation
                  supervisor = 1;                                                  // malware activation
              state = STATE_FETCH;
            end

            OPCODE_HLT: begin
              state = STATE_HALT;
            end

            default: begin
              error = 1;
              state = STATE_HALT;
            end
            
          endcase
                  
        end
      endcase
    end
  
    always@(posedge Clock) begin
      case(PC)
        6'h10: mem = {OPCODE_NOP, 4'h0 };  //
        6'h11: mem = {OPCODE_SET, 4'h1 };  //   legal out
        6'h12: mem = {OPCODE_SVC, 4'h0 };  //                           supervisor led on     
        6'h13: mem = {OPCODE_SET, 4'h2 };  //
        6'h14: mem = {OPCODE_SVC, 4'h0 };  //                           supervisor led on     
        6'h15: mem = {OPCODE_SET, 4'h4 };  //
        6'h16: mem = {OPCODE_SVC, 4'h0 };  //                           supervisor led on     
        6'h17: mem = {OPCODE_SET, 4'h8 };  //   failed out
        6'h18: mem = {OPCODE_OUT, 4'h0 };  //                           error led on
        6'h19: mem = {OPCODE_SVC, 4'h0 };  //                           supervisor led on
        6'h1A: mem = {OPCODE_SET, 4'hF };  //   
        6'h1B: mem = {OPCODE_DEC, 4'h0 };  //   troyan activation
        6'h1C: mem = {OPCODE_NOP, 4'h0 };  //   troyan activation
        6'h1D: mem = {OPCODE_JNZ, 4'h2 };  //   troyan activation       supervisor led on
        6'h1E: mem = {OPCODE_SET, 4'h1 };  //   exploitation
        6'h1F: mem = {OPCODE_OUT, 4'h0 };  //   exploitation
        6'h20: mem = {OPCODE_SET, 4'h2 };  //   exploitation
        6'h21: mem = {OPCODE_OUT, 4'h0 };  //   exploitation
        6'h22: mem = {OPCODE_SET, 4'h4 };  //   exploitation
        6'h23: mem = {OPCODE_OUT, 4'h0 };  //   exploitation
        6'h24: mem = {OPCODE_SET, 4'h8 };  //   exploitation
        6'h25: mem = {OPCODE_OUT, 4'h0 };  //   exploitation
        6'h26: mem = {OPCODE_SET, 4'h4 };  //   exploitation
        6'h27: mem = {OPCODE_OUT, 4'h0 };  //   exploitation
        6'h28: mem = {OPCODE_SET, 4'h2 };  //   exploitation
        6'h29: mem = {OPCODE_OUT, 4'h0 };  //   exploitation
        6'h2A: mem = {OPCODE_SET, 4'h1 };  //   exploitation
        6'h2B: mem = {OPCODE_OUT, 4'h0 };  //   exploitation
        6'h2C: mem = {OPCODE_NOP, 4'h0 };  //
        6'h2D: mem = {OPCODE_HLT, 4'h0 };  //
        6'h2E: mem = {OPCODE_OUT, 4'h0 };  //   svc                     gpio change
        6'h2F: mem = {OPCODE_RET, 4'h0 };  //
        default: mem = {OPCODE_HLT, 4'h0 };
      endcase
    end    

endmodule
