module board(
  input Clock,
  input reset_button,
  input step_button,
  input run_switch,
  input fast_switch,
  input malware_switch,                                          // malware enable
  input malware_input,                                           // malware manual activation
  output [7:0] SEG,
  output [7:0] DIGIT,
  
  output humanClock_led,
  output run_led,
  output supervisor_led,
  output error_led,

  output FETCH_led,
  output DECODE_led,
  output HALT_led,
  
  output NOP_led,
  output SET_led,
  output DEC_led,
  output SVC_led,
  output RET_led,
  output JNZ_led,
  output OUT_led,
  
  output malware_activation_led,                                    // malware monitoring
  output malware_activation_signal_out,                             // malware activation
  input  malware_activation_signal_in,                              // malware activation

  output [3:0] pmod_gpio

);

wire reset;
wire step;
wire run;
wire fast;

wire humanClock;

assign humanClock_led = humanClock;
assign run_led        = run;
assign supervisor_led = cpu.supervisor;
assign error_led      = cpu.error;

assign FETCH_led      = ( cpu.state == cpu.STATE_FETCH);
assign DECODE_led     = ( cpu.state == cpu.STATE_DECODE);
assign HALT_led       = ( cpu.state == cpu.STATE_HALT);
 
assign RET_led = ( cpu.opcode == cpu.OPCODE_RET ); 
assign JNZ_led = ( cpu.opcode == cpu.OPCODE_JNZ );
assign SET_led = ( cpu.opcode == cpu.OPCODE_SET );  
assign OUT_led = ( cpu.opcode == cpu.OPCODE_OUT );
assign SVC_led = ( cpu.opcode == cpu.OPCODE_SVC ); 
assign DEC_led = ( cpu.opcode == cpu.OPCODE_DEC );
assign NOP_led = ( cpu.opcode == cpu.OPCODE_NOP );

assign malware_activation_led = cpu.opcode[3];                             // malware monitoring
assign malware_activation_signal_out = cpu.opcode[3] ? 1 : 1'bz;           // malware activation


debouncer step_debouncer(.CLK(Clock),
  .switch_input(step_button),
  .state(step)
);

debouncer reset_debouncer(.CLK(Clock),
  .switch_input(reset_button),
  .state(reset)
);

debouncer run_debouncer(.CLK(Clock),
  .switch_input(run_switch),
  .state(run)
);

debouncer fast_debouncer(.CLK(Clock),
  .switch_input(fast_switch),
  .state(fast)
);

counter counter(
   .CLK(Clock),
   .reset(reset),
   .enable(run),
   .step(step),
   .fast(fast),
   .humanClock(humanClock)
);


cpu cpu(
  .Clock(humanClock),
  .reset(reset),
  .gpio(pmod_gpio)
);

display_7_seg display(.CLK (Clock),
  .number_in(
    {
     2'b00,cpu.PC,
     4'b0000,
     cpu.A[3:0],
     4'b0000,
     cpu.opcode,
     4'b0000,
     cpu.opdata
    }
  ),
  .SEG (SEG),
  .DIGIT (DIGIT)
);

endmodule
